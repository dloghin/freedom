module DecodePosit( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [31:0] io_i_bits, // @[:@6.4]
  output        io_o_posit_sign, // @[:@6.4]
  output        io_o_posit_special_number, // @[:@6.4]
  output [31:0] io_o_posit_regime, // @[:@6.4]
  output [31:0] io_o_posit_exponent, // @[:@6.4]
  output [31:0] io_o_posit_fraction, // @[:@6.4]
  output [4:0]  io_o_posit_regime_size, // @[:@6.4]
  output [4:0]  io_o_posit_exponent_size, // @[:@6.4]
  output [4:0]  io_o_posit_fraction_size, // @[:@6.4]
  output [4:0]  io_o_posit_max_exponent_size // @[:@6.4]
);
  wire  _T_14; // @[POSIT.scala 47:50:@9.4]
  wire  _T_17; // @[POSIT.scala 48:50:@11.4]
  wire [30:0] _T_25; // @[POSIT.scala 71:37:@19.4]
  wire [30:0] _T_26; // @[POSIT.scala 71:27:@20.4]
  wire [31:0] _T_28; // @[POSIT.scala 71:50:@21.4]
  wire [30:0] _T_29; // @[POSIT.scala 71:50:@22.4]
  wire [30:0] bits_to_decode; // @[POSIT.scala 70:26:@24.4]
  wire  _T_33; // @[POSIT.scala 80:51:@27.4]
  wire [30:0] _T_34; // @[POSIT.scala 81:61:@28.4]
  wire [15:0] _T_35; // @[Bitwise.scala 109:18:@29.4]
  wire [7:0] _T_40; // @[Bitwise.scala 103:21:@32.4]
  wire [15:0] _T_41; // @[Bitwise.scala 103:31:@33.4]
  wire [7:0] _T_42; // @[Bitwise.scala 103:46:@34.4]
  wire [15:0] _GEN_0; // @[Bitwise.scala 103:65:@35.4]
  wire [15:0] _T_43; // @[Bitwise.scala 103:65:@35.4]
  wire [15:0] _T_45; // @[Bitwise.scala 103:75:@37.4]
  wire [15:0] _T_46; // @[Bitwise.scala 103:39:@38.4]
  wire [11:0] _T_50; // @[Bitwise.scala 103:21:@42.4]
  wire [15:0] _GEN_1; // @[Bitwise.scala 103:31:@43.4]
  wire [15:0] _T_51; // @[Bitwise.scala 103:31:@43.4]
  wire [11:0] _T_52; // @[Bitwise.scala 103:46:@44.4]
  wire [15:0] _GEN_2; // @[Bitwise.scala 103:65:@45.4]
  wire [15:0] _T_53; // @[Bitwise.scala 103:65:@45.4]
  wire [15:0] _T_55; // @[Bitwise.scala 103:75:@47.4]
  wire [15:0] _T_56; // @[Bitwise.scala 103:39:@48.4]
  wire [13:0] _T_60; // @[Bitwise.scala 103:21:@52.4]
  wire [15:0] _GEN_3; // @[Bitwise.scala 103:31:@53.4]
  wire [15:0] _T_61; // @[Bitwise.scala 103:31:@53.4]
  wire [13:0] _T_62; // @[Bitwise.scala 103:46:@54.4]
  wire [15:0] _GEN_4; // @[Bitwise.scala 103:65:@55.4]
  wire [15:0] _T_63; // @[Bitwise.scala 103:65:@55.4]
  wire [15:0] _T_65; // @[Bitwise.scala 103:75:@57.4]
  wire [15:0] _T_66; // @[Bitwise.scala 103:39:@58.4]
  wire [14:0] _T_70; // @[Bitwise.scala 103:21:@62.4]
  wire [15:0] _GEN_5; // @[Bitwise.scala 103:31:@63.4]
  wire [15:0] _T_71; // @[Bitwise.scala 103:31:@63.4]
  wire [14:0] _T_72; // @[Bitwise.scala 103:46:@64.4]
  wire [15:0] _GEN_6; // @[Bitwise.scala 103:65:@65.4]
  wire [15:0] _T_73; // @[Bitwise.scala 103:65:@65.4]
  wire [15:0] _T_75; // @[Bitwise.scala 103:75:@67.4]
  wire [15:0] _T_76; // @[Bitwise.scala 103:39:@68.4]
  wire [14:0] _T_77; // @[Bitwise.scala 109:44:@69.4]
  wire [7:0] _T_78; // @[Bitwise.scala 109:18:@70.4]
  wire [3:0] _T_83; // @[Bitwise.scala 103:21:@73.4]
  wire [7:0] _T_84; // @[Bitwise.scala 103:31:@74.4]
  wire [3:0] _T_85; // @[Bitwise.scala 103:46:@75.4]
  wire [7:0] _GEN_7; // @[Bitwise.scala 103:65:@76.4]
  wire [7:0] _T_86; // @[Bitwise.scala 103:65:@76.4]
  wire [7:0] _T_88; // @[Bitwise.scala 103:75:@78.4]
  wire [7:0] _T_89; // @[Bitwise.scala 103:39:@79.4]
  wire [5:0] _T_93; // @[Bitwise.scala 103:21:@83.4]
  wire [7:0] _GEN_8; // @[Bitwise.scala 103:31:@84.4]
  wire [7:0] _T_94; // @[Bitwise.scala 103:31:@84.4]
  wire [5:0] _T_95; // @[Bitwise.scala 103:46:@85.4]
  wire [7:0] _GEN_9; // @[Bitwise.scala 103:65:@86.4]
  wire [7:0] _T_96; // @[Bitwise.scala 103:65:@86.4]
  wire [7:0] _T_98; // @[Bitwise.scala 103:75:@88.4]
  wire [7:0] _T_99; // @[Bitwise.scala 103:39:@89.4]
  wire [6:0] _T_103; // @[Bitwise.scala 103:21:@93.4]
  wire [7:0] _GEN_10; // @[Bitwise.scala 103:31:@94.4]
  wire [7:0] _T_104; // @[Bitwise.scala 103:31:@94.4]
  wire [6:0] _T_105; // @[Bitwise.scala 103:46:@95.4]
  wire [7:0] _GEN_11; // @[Bitwise.scala 103:65:@96.4]
  wire [7:0] _T_106; // @[Bitwise.scala 103:65:@96.4]
  wire [7:0] _T_108; // @[Bitwise.scala 103:75:@98.4]
  wire [7:0] _T_109; // @[Bitwise.scala 103:39:@99.4]
  wire [6:0] _T_110; // @[Bitwise.scala 109:44:@100.4]
  wire [3:0] _T_111; // @[Bitwise.scala 109:18:@101.4]
  wire [1:0] _T_112; // @[Bitwise.scala 109:18:@102.4]
  wire  _T_113; // @[Bitwise.scala 109:18:@103.4]
  wire  _T_114; // @[Bitwise.scala 109:44:@104.4]
  wire [1:0] _T_116; // @[Bitwise.scala 109:44:@106.4]
  wire  _T_117; // @[Bitwise.scala 109:18:@107.4]
  wire  _T_118; // @[Bitwise.scala 109:44:@108.4]
  wire [2:0] _T_121; // @[Bitwise.scala 109:44:@111.4]
  wire [1:0] _T_122; // @[Bitwise.scala 109:18:@112.4]
  wire  _T_123; // @[Bitwise.scala 109:18:@113.4]
  wire  _T_124; // @[Bitwise.scala 109:44:@114.4]
  wire  _T_126; // @[Bitwise.scala 109:44:@116.4]
  wire [30:0] _T_130; // @[Cat.scala 30:58:@120.4]
  wire  _T_131; // @[OneHot.scala 39:40:@121.4]
  wire  _T_132; // @[OneHot.scala 39:40:@122.4]
  wire  _T_133; // @[OneHot.scala 39:40:@123.4]
  wire  _T_134; // @[OneHot.scala 39:40:@124.4]
  wire  _T_135; // @[OneHot.scala 39:40:@125.4]
  wire  _T_136; // @[OneHot.scala 39:40:@126.4]
  wire  _T_137; // @[OneHot.scala 39:40:@127.4]
  wire  _T_138; // @[OneHot.scala 39:40:@128.4]
  wire  _T_139; // @[OneHot.scala 39:40:@129.4]
  wire  _T_140; // @[OneHot.scala 39:40:@130.4]
  wire  _T_141; // @[OneHot.scala 39:40:@131.4]
  wire  _T_142; // @[OneHot.scala 39:40:@132.4]
  wire  _T_143; // @[OneHot.scala 39:40:@133.4]
  wire  _T_144; // @[OneHot.scala 39:40:@134.4]
  wire  _T_145; // @[OneHot.scala 39:40:@135.4]
  wire  _T_146; // @[OneHot.scala 39:40:@136.4]
  wire  _T_147; // @[OneHot.scala 39:40:@137.4]
  wire  _T_148; // @[OneHot.scala 39:40:@138.4]
  wire  _T_149; // @[OneHot.scala 39:40:@139.4]
  wire  _T_150; // @[OneHot.scala 39:40:@140.4]
  wire  _T_151; // @[OneHot.scala 39:40:@141.4]
  wire  _T_152; // @[OneHot.scala 39:40:@142.4]
  wire  _T_153; // @[OneHot.scala 39:40:@143.4]
  wire  _T_154; // @[OneHot.scala 39:40:@144.4]
  wire  _T_155; // @[OneHot.scala 39:40:@145.4]
  wire  _T_156; // @[OneHot.scala 39:40:@146.4]
  wire  _T_157; // @[OneHot.scala 39:40:@147.4]
  wire  _T_158; // @[OneHot.scala 39:40:@148.4]
  wire  _T_159; // @[OneHot.scala 39:40:@149.4]
  wire  _T_160; // @[OneHot.scala 39:40:@150.4]
  wire [4:0] _T_193; // @[Mux.scala 31:69:@152.4]
  wire [4:0] _T_194; // @[Mux.scala 31:69:@153.4]
  wire [4:0] _T_195; // @[Mux.scala 31:69:@154.4]
  wire [4:0] _T_196; // @[Mux.scala 31:69:@155.4]
  wire [4:0] _T_197; // @[Mux.scala 31:69:@156.4]
  wire [4:0] _T_198; // @[Mux.scala 31:69:@157.4]
  wire [4:0] _T_199; // @[Mux.scala 31:69:@158.4]
  wire [4:0] _T_200; // @[Mux.scala 31:69:@159.4]
  wire [4:0] _T_201; // @[Mux.scala 31:69:@160.4]
  wire [4:0] _T_202; // @[Mux.scala 31:69:@161.4]
  wire [4:0] _T_203; // @[Mux.scala 31:69:@162.4]
  wire [4:0] _T_204; // @[Mux.scala 31:69:@163.4]
  wire [4:0] _T_205; // @[Mux.scala 31:69:@164.4]
  wire [4:0] _T_206; // @[Mux.scala 31:69:@165.4]
  wire [4:0] _T_207; // @[Mux.scala 31:69:@166.4]
  wire [4:0] _T_208; // @[Mux.scala 31:69:@167.4]
  wire [4:0] _T_209; // @[Mux.scala 31:69:@168.4]
  wire [4:0] _T_210; // @[Mux.scala 31:69:@169.4]
  wire [4:0] _T_211; // @[Mux.scala 31:69:@170.4]
  wire [4:0] _T_212; // @[Mux.scala 31:69:@171.4]
  wire [4:0] _T_213; // @[Mux.scala 31:69:@172.4]
  wire [4:0] _T_214; // @[Mux.scala 31:69:@173.4]
  wire [4:0] _T_215; // @[Mux.scala 31:69:@174.4]
  wire [4:0] _T_216; // @[Mux.scala 31:69:@175.4]
  wire [4:0] _T_217; // @[Mux.scala 31:69:@176.4]
  wire [4:0] _T_218; // @[Mux.scala 31:69:@177.4]
  wire [4:0] _T_219; // @[Mux.scala 31:69:@178.4]
  wire [4:0] _T_220; // @[Mux.scala 31:69:@179.4]
  wire [4:0] _T_221; // @[Mux.scala 31:69:@180.4]
  wire [4:0] _T_222; // @[Mux.scala 31:69:@181.4]
  wire [15:0] _T_223; // @[Bitwise.scala 109:18:@182.4]
  wire [7:0] _T_228; // @[Bitwise.scala 103:21:@185.4]
  wire [15:0] _T_229; // @[Bitwise.scala 103:31:@186.4]
  wire [7:0] _T_230; // @[Bitwise.scala 103:46:@187.4]
  wire [15:0] _GEN_12; // @[Bitwise.scala 103:65:@188.4]
  wire [15:0] _T_231; // @[Bitwise.scala 103:65:@188.4]
  wire [15:0] _T_233; // @[Bitwise.scala 103:75:@190.4]
  wire [15:0] _T_234; // @[Bitwise.scala 103:39:@191.4]
  wire [11:0] _T_238; // @[Bitwise.scala 103:21:@195.4]
  wire [15:0] _GEN_13; // @[Bitwise.scala 103:31:@196.4]
  wire [15:0] _T_239; // @[Bitwise.scala 103:31:@196.4]
  wire [11:0] _T_240; // @[Bitwise.scala 103:46:@197.4]
  wire [15:0] _GEN_14; // @[Bitwise.scala 103:65:@198.4]
  wire [15:0] _T_241; // @[Bitwise.scala 103:65:@198.4]
  wire [15:0] _T_243; // @[Bitwise.scala 103:75:@200.4]
  wire [15:0] _T_244; // @[Bitwise.scala 103:39:@201.4]
  wire [13:0] _T_248; // @[Bitwise.scala 103:21:@205.4]
  wire [15:0] _GEN_15; // @[Bitwise.scala 103:31:@206.4]
  wire [15:0] _T_249; // @[Bitwise.scala 103:31:@206.4]
  wire [13:0] _T_250; // @[Bitwise.scala 103:46:@207.4]
  wire [15:0] _GEN_16; // @[Bitwise.scala 103:65:@208.4]
  wire [15:0] _T_251; // @[Bitwise.scala 103:65:@208.4]
  wire [15:0] _T_253; // @[Bitwise.scala 103:75:@210.4]
  wire [15:0] _T_254; // @[Bitwise.scala 103:39:@211.4]
  wire [14:0] _T_258; // @[Bitwise.scala 103:21:@215.4]
  wire [15:0] _GEN_17; // @[Bitwise.scala 103:31:@216.4]
  wire [15:0] _T_259; // @[Bitwise.scala 103:31:@216.4]
  wire [14:0] _T_260; // @[Bitwise.scala 103:46:@217.4]
  wire [15:0] _GEN_18; // @[Bitwise.scala 103:65:@218.4]
  wire [15:0] _T_261; // @[Bitwise.scala 103:65:@218.4]
  wire [15:0] _T_263; // @[Bitwise.scala 103:75:@220.4]
  wire [15:0] _T_264; // @[Bitwise.scala 103:39:@221.4]
  wire [14:0] _T_265; // @[Bitwise.scala 109:44:@222.4]
  wire [7:0] _T_266; // @[Bitwise.scala 109:18:@223.4]
  wire [3:0] _T_271; // @[Bitwise.scala 103:21:@226.4]
  wire [7:0] _T_272; // @[Bitwise.scala 103:31:@227.4]
  wire [3:0] _T_273; // @[Bitwise.scala 103:46:@228.4]
  wire [7:0] _GEN_19; // @[Bitwise.scala 103:65:@229.4]
  wire [7:0] _T_274; // @[Bitwise.scala 103:65:@229.4]
  wire [7:0] _T_276; // @[Bitwise.scala 103:75:@231.4]
  wire [7:0] _T_277; // @[Bitwise.scala 103:39:@232.4]
  wire [5:0] _T_281; // @[Bitwise.scala 103:21:@236.4]
  wire [7:0] _GEN_20; // @[Bitwise.scala 103:31:@237.4]
  wire [7:0] _T_282; // @[Bitwise.scala 103:31:@237.4]
  wire [5:0] _T_283; // @[Bitwise.scala 103:46:@238.4]
  wire [7:0] _GEN_21; // @[Bitwise.scala 103:65:@239.4]
  wire [7:0] _T_284; // @[Bitwise.scala 103:65:@239.4]
  wire [7:0] _T_286; // @[Bitwise.scala 103:75:@241.4]
  wire [7:0] _T_287; // @[Bitwise.scala 103:39:@242.4]
  wire [6:0] _T_291; // @[Bitwise.scala 103:21:@246.4]
  wire [7:0] _GEN_22; // @[Bitwise.scala 103:31:@247.4]
  wire [7:0] _T_292; // @[Bitwise.scala 103:31:@247.4]
  wire [6:0] _T_293; // @[Bitwise.scala 103:46:@248.4]
  wire [7:0] _GEN_23; // @[Bitwise.scala 103:65:@249.4]
  wire [7:0] _T_294; // @[Bitwise.scala 103:65:@249.4]
  wire [7:0] _T_296; // @[Bitwise.scala 103:75:@251.4]
  wire [7:0] _T_297; // @[Bitwise.scala 103:39:@252.4]
  wire [6:0] _T_298; // @[Bitwise.scala 109:44:@253.4]
  wire [3:0] _T_299; // @[Bitwise.scala 109:18:@254.4]
  wire [1:0] _T_300; // @[Bitwise.scala 109:18:@255.4]
  wire  _T_301; // @[Bitwise.scala 109:18:@256.4]
  wire  _T_302; // @[Bitwise.scala 109:44:@257.4]
  wire [1:0] _T_304; // @[Bitwise.scala 109:44:@259.4]
  wire  _T_305; // @[Bitwise.scala 109:18:@260.4]
  wire  _T_306; // @[Bitwise.scala 109:44:@261.4]
  wire [2:0] _T_309; // @[Bitwise.scala 109:44:@264.4]
  wire [1:0] _T_310; // @[Bitwise.scala 109:18:@265.4]
  wire  _T_311; // @[Bitwise.scala 109:18:@266.4]
  wire  _T_312; // @[Bitwise.scala 109:44:@267.4]
  wire  _T_314; // @[Bitwise.scala 109:44:@269.4]
  wire [30:0] _T_318; // @[Cat.scala 30:58:@273.4]
  wire  _T_319; // @[OneHot.scala 39:40:@274.4]
  wire  _T_320; // @[OneHot.scala 39:40:@275.4]
  wire  _T_321; // @[OneHot.scala 39:40:@276.4]
  wire  _T_322; // @[OneHot.scala 39:40:@277.4]
  wire  _T_323; // @[OneHot.scala 39:40:@278.4]
  wire  _T_324; // @[OneHot.scala 39:40:@279.4]
  wire  _T_325; // @[OneHot.scala 39:40:@280.4]
  wire  _T_326; // @[OneHot.scala 39:40:@281.4]
  wire  _T_327; // @[OneHot.scala 39:40:@282.4]
  wire  _T_328; // @[OneHot.scala 39:40:@283.4]
  wire  _T_329; // @[OneHot.scala 39:40:@284.4]
  wire  _T_330; // @[OneHot.scala 39:40:@285.4]
  wire  _T_331; // @[OneHot.scala 39:40:@286.4]
  wire  _T_332; // @[OneHot.scala 39:40:@287.4]
  wire  _T_333; // @[OneHot.scala 39:40:@288.4]
  wire  _T_334; // @[OneHot.scala 39:40:@289.4]
  wire  _T_335; // @[OneHot.scala 39:40:@290.4]
  wire  _T_336; // @[OneHot.scala 39:40:@291.4]
  wire  _T_337; // @[OneHot.scala 39:40:@292.4]
  wire  _T_338; // @[OneHot.scala 39:40:@293.4]
  wire  _T_339; // @[OneHot.scala 39:40:@294.4]
  wire  _T_340; // @[OneHot.scala 39:40:@295.4]
  wire  _T_341; // @[OneHot.scala 39:40:@296.4]
  wire  _T_342; // @[OneHot.scala 39:40:@297.4]
  wire  _T_343; // @[OneHot.scala 39:40:@298.4]
  wire  _T_344; // @[OneHot.scala 39:40:@299.4]
  wire  _T_345; // @[OneHot.scala 39:40:@300.4]
  wire  _T_346; // @[OneHot.scala 39:40:@301.4]
  wire  _T_347; // @[OneHot.scala 39:40:@302.4]
  wire  _T_348; // @[OneHot.scala 39:40:@303.4]
  wire [4:0] _T_381; // @[Mux.scala 31:69:@305.4]
  wire [4:0] _T_382; // @[Mux.scala 31:69:@306.4]
  wire [4:0] _T_383; // @[Mux.scala 31:69:@307.4]
  wire [4:0] _T_384; // @[Mux.scala 31:69:@308.4]
  wire [4:0] _T_385; // @[Mux.scala 31:69:@309.4]
  wire [4:0] _T_386; // @[Mux.scala 31:69:@310.4]
  wire [4:0] _T_387; // @[Mux.scala 31:69:@311.4]
  wire [4:0] _T_388; // @[Mux.scala 31:69:@312.4]
  wire [4:0] _T_389; // @[Mux.scala 31:69:@313.4]
  wire [4:0] _T_390; // @[Mux.scala 31:69:@314.4]
  wire [4:0] _T_391; // @[Mux.scala 31:69:@315.4]
  wire [4:0] _T_392; // @[Mux.scala 31:69:@316.4]
  wire [4:0] _T_393; // @[Mux.scala 31:69:@317.4]
  wire [4:0] _T_394; // @[Mux.scala 31:69:@318.4]
  wire [4:0] _T_395; // @[Mux.scala 31:69:@319.4]
  wire [4:0] _T_396; // @[Mux.scala 31:69:@320.4]
  wire [4:0] _T_397; // @[Mux.scala 31:69:@321.4]
  wire [4:0] _T_398; // @[Mux.scala 31:69:@322.4]
  wire [4:0] _T_399; // @[Mux.scala 31:69:@323.4]
  wire [4:0] _T_400; // @[Mux.scala 31:69:@324.4]
  wire [4:0] _T_401; // @[Mux.scala 31:69:@325.4]
  wire [4:0] _T_402; // @[Mux.scala 31:69:@326.4]
  wire [4:0] _T_403; // @[Mux.scala 31:69:@327.4]
  wire [4:0] _T_404; // @[Mux.scala 31:69:@328.4]
  wire [4:0] _T_405; // @[Mux.scala 31:69:@329.4]
  wire [4:0] _T_406; // @[Mux.scala 31:69:@330.4]
  wire [4:0] _T_407; // @[Mux.scala 31:69:@331.4]
  wire [4:0] _T_408; // @[Mux.scala 31:69:@332.4]
  wire [4:0] _T_409; // @[Mux.scala 31:69:@333.4]
  wire [4:0] _T_410; // @[Mux.scala 31:69:@334.4]
  wire [4:0] number_of_same_bit_value; // @[POSIT.scala 80:36:@335.4]
  wire  _T_413; // @[POSIT.scala 98:47:@338.4]
  wire  _T_417; // @[POSIT.scala 98:84:@340.4]
  wire  _T_418; // @[POSIT.scala 98:57:@341.4]
  wire [5:0] _T_419; // @[POSIT.scala 99:58:@342.4]
  wire [6:0] _T_422; // @[POSIT.scala 100:63:@344.4]
  wire [5:0] _T_423; // @[POSIT.scala 100:63:@345.4]
  wire [5:0] _T_424; // @[POSIT.scala 100:63:@346.4]
  wire [5:0] _T_425; // @[POSIT.scala 98:32:@347.4]
  wire  _T_428; // @[POSIT.scala 101:51:@349.4]
  wire  _T_431; // @[POSIT.scala 101:58:@351.4]
  wire [6:0] _T_434; // @[POSIT.scala 102:30:@353.4]
  wire [5:0] _T_435; // @[POSIT.scala 102:30:@354.4]
  wire [5:0] _T_436; // @[POSIT.scala 102:30:@355.4]
  wire [6:0] _T_438; // @[POSIT.scala 102:61:@356.4]
  wire [5:0] _T_439; // @[POSIT.scala 102:61:@357.4]
  wire [5:0] _T_440; // @[POSIT.scala 102:61:@358.4]
  wire [5:0] _T_446; // @[POSIT.scala 101:33:@363.4]
  wire [5:0] _T_447; // @[POSIT.scala 97:29:@364.4]
  wire [5:0] _T_449; // @[POSIT.scala 108:56:@366.4]
  wire [7:0] _T_454; // @[POSIT.scala 116:37:@370.4]
  wire [6:0] _T_455; // @[POSIT.scala 116:37:@371.4]
  wire [6:0] _T_456; // @[POSIT.scala 116:37:@372.4]
  wire [5:0] _T_457; // @[POSIT.scala 116:68:@373.4]
  wire [6:0] _GEN_24; // @[POSIT.scala 116:43:@374.4]
  wire [7:0] _T_458; // @[POSIT.scala 116:43:@374.4]
  wire [6:0] _T_459; // @[POSIT.scala 116:43:@375.4]
  wire [6:0] _T_460; // @[POSIT.scala 116:43:@376.4]
  wire [5:0] _T_461; // @[POSIT.scala 116:104:@377.4]
  wire [6:0] _GEN_25; // @[POSIT.scala 116:73:@378.4]
  wire [7:0] _T_462; // @[POSIT.scala 116:73:@378.4]
  wire [6:0] _T_463; // @[POSIT.scala 116:73:@379.4]
  wire [6:0] _T_464; // @[POSIT.scala 116:73:@380.4]
  wire [5:0] _GEN_26; // @[POSIT.scala 115:37:@369.4 POSIT.scala 116:27:@381.4]
  wire [5:0] posible_fraction_size; // @[POSIT.scala 115:37:@369.4 POSIT.scala 116:27:@381.4]
  wire  _T_466; // @[POSIT.scala 117:59:@382.4]
  wire [6:0] _T_470; // @[POSIT.scala 119:44:@383.4]
  wire [6:0] _T_471; // @[POSIT.scala 119:44:@384.4]
  wire [5:0] _T_472; // @[POSIT.scala 119:44:@385.4]
  wire [5:0] _GEN_27; // @[POSIT.scala 119:50:@386.4]
  wire [6:0] _T_473; // @[POSIT.scala 119:50:@386.4]
  wire [6:0] _T_474; // @[POSIT.scala 119:50:@387.4]
  wire [5:0] _T_475; // @[POSIT.scala 119:50:@388.4]
  wire [5:0] _GEN_28; // @[POSIT.scala 119:75:@389.4]
  wire [6:0] _T_476; // @[POSIT.scala 119:75:@389.4]
  wire [6:0] _T_477; // @[POSIT.scala 119:75:@390.4]
  wire [5:0] _T_478; // @[POSIT.scala 119:75:@391.4]
  wire [5:0] _T_479; // @[POSIT.scala 117:36:@392.4]
  wire  _T_481; // @[POSIT.scala 124:57:@394.4]
  wire [5:0] _GEN_29; // @[POSIT.scala 126:65:@396.4]
  wire [6:0] _T_489; // @[POSIT.scala 126:65:@396.4]
  wire [6:0] _T_490; // @[POSIT.scala 126:65:@397.4]
  wire [5:0] _T_491; // @[POSIT.scala 126:65:@398.4]
  wire [31:0] _T_492; // @[POSIT.scala 126:55:@399.4]
  wire [31:0] _GEN_30; // @[POSIT.scala 126:92:@400.4]
  wire [31:0] _T_493; // @[POSIT.scala 126:92:@400.4]
  wire [5:0] _GEN_32; // @[POSIT.scala 131:39:@403.4 POSIT.scala 132:29:@411.4]
  wire [5:0] posible_exponent_size_1; // @[POSIT.scala 131:39:@403.4 POSIT.scala 132:29:@411.4]
  wire  _T_507; // @[POSIT.scala 134:60:@414.4]
  wire [5:0] posible_exponent_size_2; // @[POSIT.scala 134:35:@416.4]
  wire  _T_511; // @[POSIT.scala 137:61:@418.4]
  wire [5:0] _T_513; // @[POSIT.scala 139:61:@419.4]
  wire [5:0] _T_514; // @[POSIT.scala 137:36:@420.4]
  wire  _T_516; // @[POSIT.scala 146:57:@422.4]
  wire [30:0] _T_518; // @[POSIT.scala 148:48:@423.4]
  wire [5:0] _GEN_33; // @[POSIT.scala 149:64:@425.4]
  wire [6:0] _T_525; // @[POSIT.scala 149:64:@425.4]
  wire [6:0] _T_526; // @[POSIT.scala 149:64:@426.4]
  wire [5:0] _T_527; // @[POSIT.scala 149:64:@427.4]
  wire [31:0] _T_528; // @[POSIT.scala 149:53:@428.4]
  wire [31:0] _GEN_34; // @[POSIT.scala 148:79:@429.4]
  wire [31:0] _T_529; // @[POSIT.scala 148:79:@429.4]
  assign _T_14 = io_i_bits == 32'h0; // @[POSIT.scala 47:50:@9.4]
  assign _T_17 = io_i_bits == 32'h80000000; // @[POSIT.scala 48:50:@11.4]
  assign _T_25 = io_i_bits[30:0]; // @[POSIT.scala 71:37:@19.4]
  assign _T_26 = ~ _T_25; // @[POSIT.scala 71:27:@20.4]
  assign _T_28 = _T_26 + 31'h1; // @[POSIT.scala 71:50:@21.4]
  assign _T_29 = _T_26 + 31'h1; // @[POSIT.scala 71:50:@22.4]
  assign bits_to_decode = io_o_posit_sign ? _T_29 : _T_25; // @[POSIT.scala 70:26:@24.4]
  assign _T_33 = bits_to_decode[30]; // @[POSIT.scala 80:51:@27.4]
  assign _T_34 = ~ bits_to_decode; // @[POSIT.scala 81:61:@28.4]
  assign _T_35 = _T_34[15:0]; // @[Bitwise.scala 109:18:@29.4]
  assign _T_40 = _T_35[15:8]; // @[Bitwise.scala 103:21:@32.4]
  assign _T_41 = {{8'd0}, _T_40}; // @[Bitwise.scala 103:31:@33.4]
  assign _T_42 = _T_35[7:0]; // @[Bitwise.scala 103:46:@34.4]
  assign _GEN_0 = {{8'd0}, _T_42}; // @[Bitwise.scala 103:65:@35.4]
  assign _T_43 = _GEN_0 << 8; // @[Bitwise.scala 103:65:@35.4]
  assign _T_45 = _T_43 & 16'hff00; // @[Bitwise.scala 103:75:@37.4]
  assign _T_46 = _T_41 | _T_45; // @[Bitwise.scala 103:39:@38.4]
  assign _T_50 = _T_46[15:4]; // @[Bitwise.scala 103:21:@42.4]
  assign _GEN_1 = {{4'd0}, _T_50}; // @[Bitwise.scala 103:31:@43.4]
  assign _T_51 = _GEN_1 & 16'hf0f; // @[Bitwise.scala 103:31:@43.4]
  assign _T_52 = _T_46[11:0]; // @[Bitwise.scala 103:46:@44.4]
  assign _GEN_2 = {{4'd0}, _T_52}; // @[Bitwise.scala 103:65:@45.4]
  assign _T_53 = _GEN_2 << 4; // @[Bitwise.scala 103:65:@45.4]
  assign _T_55 = _T_53 & 16'hf0f0; // @[Bitwise.scala 103:75:@47.4]
  assign _T_56 = _T_51 | _T_55; // @[Bitwise.scala 103:39:@48.4]
  assign _T_60 = _T_56[15:2]; // @[Bitwise.scala 103:21:@52.4]
  assign _GEN_3 = {{2'd0}, _T_60}; // @[Bitwise.scala 103:31:@53.4]
  assign _T_61 = _GEN_3 & 16'h3333; // @[Bitwise.scala 103:31:@53.4]
  assign _T_62 = _T_56[13:0]; // @[Bitwise.scala 103:46:@54.4]
  assign _GEN_4 = {{2'd0}, _T_62}; // @[Bitwise.scala 103:65:@55.4]
  assign _T_63 = _GEN_4 << 2; // @[Bitwise.scala 103:65:@55.4]
  assign _T_65 = _T_63 & 16'hcccc; // @[Bitwise.scala 103:75:@57.4]
  assign _T_66 = _T_61 | _T_65; // @[Bitwise.scala 103:39:@58.4]
  assign _T_70 = _T_66[15:1]; // @[Bitwise.scala 103:21:@62.4]
  assign _GEN_5 = {{1'd0}, _T_70}; // @[Bitwise.scala 103:31:@63.4]
  assign _T_71 = _GEN_5 & 16'h5555; // @[Bitwise.scala 103:31:@63.4]
  assign _T_72 = _T_66[14:0]; // @[Bitwise.scala 103:46:@64.4]
  assign _GEN_6 = {{1'd0}, _T_72}; // @[Bitwise.scala 103:65:@65.4]
  assign _T_73 = _GEN_6 << 1; // @[Bitwise.scala 103:65:@65.4]
  assign _T_75 = _T_73 & 16'haaaa; // @[Bitwise.scala 103:75:@67.4]
  assign _T_76 = _T_71 | _T_75; // @[Bitwise.scala 103:39:@68.4]
  assign _T_77 = _T_34[30:16]; // @[Bitwise.scala 109:44:@69.4]
  assign _T_78 = _T_77[7:0]; // @[Bitwise.scala 109:18:@70.4]
  assign _T_83 = _T_78[7:4]; // @[Bitwise.scala 103:21:@73.4]
  assign _T_84 = {{4'd0}, _T_83}; // @[Bitwise.scala 103:31:@74.4]
  assign _T_85 = _T_78[3:0]; // @[Bitwise.scala 103:46:@75.4]
  assign _GEN_7 = {{4'd0}, _T_85}; // @[Bitwise.scala 103:65:@76.4]
  assign _T_86 = _GEN_7 << 4; // @[Bitwise.scala 103:65:@76.4]
  assign _T_88 = _T_86 & 8'hf0; // @[Bitwise.scala 103:75:@78.4]
  assign _T_89 = _T_84 | _T_88; // @[Bitwise.scala 103:39:@79.4]
  assign _T_93 = _T_89[7:2]; // @[Bitwise.scala 103:21:@83.4]
  assign _GEN_8 = {{2'd0}, _T_93}; // @[Bitwise.scala 103:31:@84.4]
  assign _T_94 = _GEN_8 & 8'h33; // @[Bitwise.scala 103:31:@84.4]
  assign _T_95 = _T_89[5:0]; // @[Bitwise.scala 103:46:@85.4]
  assign _GEN_9 = {{2'd0}, _T_95}; // @[Bitwise.scala 103:65:@86.4]
  assign _T_96 = _GEN_9 << 2; // @[Bitwise.scala 103:65:@86.4]
  assign _T_98 = _T_96 & 8'hcc; // @[Bitwise.scala 103:75:@88.4]
  assign _T_99 = _T_94 | _T_98; // @[Bitwise.scala 103:39:@89.4]
  assign _T_103 = _T_99[7:1]; // @[Bitwise.scala 103:21:@93.4]
  assign _GEN_10 = {{1'd0}, _T_103}; // @[Bitwise.scala 103:31:@94.4]
  assign _T_104 = _GEN_10 & 8'h55; // @[Bitwise.scala 103:31:@94.4]
  assign _T_105 = _T_99[6:0]; // @[Bitwise.scala 103:46:@95.4]
  assign _GEN_11 = {{1'd0}, _T_105}; // @[Bitwise.scala 103:65:@96.4]
  assign _T_106 = _GEN_11 << 1; // @[Bitwise.scala 103:65:@96.4]
  assign _T_108 = _T_106 & 8'haa; // @[Bitwise.scala 103:75:@98.4]
  assign _T_109 = _T_104 | _T_108; // @[Bitwise.scala 103:39:@99.4]
  assign _T_110 = _T_77[14:8]; // @[Bitwise.scala 109:44:@100.4]
  assign _T_111 = _T_110[3:0]; // @[Bitwise.scala 109:18:@101.4]
  assign _T_112 = _T_111[1:0]; // @[Bitwise.scala 109:18:@102.4]
  assign _T_113 = _T_112[0]; // @[Bitwise.scala 109:18:@103.4]
  assign _T_114 = _T_112[1]; // @[Bitwise.scala 109:44:@104.4]
  assign _T_116 = _T_111[3:2]; // @[Bitwise.scala 109:44:@106.4]
  assign _T_117 = _T_116[0]; // @[Bitwise.scala 109:18:@107.4]
  assign _T_118 = _T_116[1]; // @[Bitwise.scala 109:44:@108.4]
  assign _T_121 = _T_110[6:4]; // @[Bitwise.scala 109:44:@111.4]
  assign _T_122 = _T_121[1:0]; // @[Bitwise.scala 109:18:@112.4]
  assign _T_123 = _T_122[0]; // @[Bitwise.scala 109:18:@113.4]
  assign _T_124 = _T_122[1]; // @[Bitwise.scala 109:44:@114.4]
  assign _T_126 = _T_121[2]; // @[Bitwise.scala 109:44:@116.4]
  assign _T_130 = {_T_76,_T_109,_T_113,_T_114,_T_117,_T_118,_T_123,_T_124,_T_126}; // @[Cat.scala 30:58:@120.4]
  assign _T_131 = _T_130[0]; // @[OneHot.scala 39:40:@121.4]
  assign _T_132 = _T_130[1]; // @[OneHot.scala 39:40:@122.4]
  assign _T_133 = _T_130[2]; // @[OneHot.scala 39:40:@123.4]
  assign _T_134 = _T_130[3]; // @[OneHot.scala 39:40:@124.4]
  assign _T_135 = _T_130[4]; // @[OneHot.scala 39:40:@125.4]
  assign _T_136 = _T_130[5]; // @[OneHot.scala 39:40:@126.4]
  assign _T_137 = _T_130[6]; // @[OneHot.scala 39:40:@127.4]
  assign _T_138 = _T_130[7]; // @[OneHot.scala 39:40:@128.4]
  assign _T_139 = _T_130[8]; // @[OneHot.scala 39:40:@129.4]
  assign _T_140 = _T_130[9]; // @[OneHot.scala 39:40:@130.4]
  assign _T_141 = _T_130[10]; // @[OneHot.scala 39:40:@131.4]
  assign _T_142 = _T_130[11]; // @[OneHot.scala 39:40:@132.4]
  assign _T_143 = _T_130[12]; // @[OneHot.scala 39:40:@133.4]
  assign _T_144 = _T_130[13]; // @[OneHot.scala 39:40:@134.4]
  assign _T_145 = _T_130[14]; // @[OneHot.scala 39:40:@135.4]
  assign _T_146 = _T_130[15]; // @[OneHot.scala 39:40:@136.4]
  assign _T_147 = _T_130[16]; // @[OneHot.scala 39:40:@137.4]
  assign _T_148 = _T_130[17]; // @[OneHot.scala 39:40:@138.4]
  assign _T_149 = _T_130[18]; // @[OneHot.scala 39:40:@139.4]
  assign _T_150 = _T_130[19]; // @[OneHot.scala 39:40:@140.4]
  assign _T_151 = _T_130[20]; // @[OneHot.scala 39:40:@141.4]
  assign _T_152 = _T_130[21]; // @[OneHot.scala 39:40:@142.4]
  assign _T_153 = _T_130[22]; // @[OneHot.scala 39:40:@143.4]
  assign _T_154 = _T_130[23]; // @[OneHot.scala 39:40:@144.4]
  assign _T_155 = _T_130[24]; // @[OneHot.scala 39:40:@145.4]
  assign _T_156 = _T_130[25]; // @[OneHot.scala 39:40:@146.4]
  assign _T_157 = _T_130[26]; // @[OneHot.scala 39:40:@147.4]
  assign _T_158 = _T_130[27]; // @[OneHot.scala 39:40:@148.4]
  assign _T_159 = _T_130[28]; // @[OneHot.scala 39:40:@149.4]
  assign _T_160 = _T_130[29]; // @[OneHot.scala 39:40:@150.4]
  assign _T_193 = _T_160 ? 5'h1d : 5'h1e; // @[Mux.scala 31:69:@152.4]
  assign _T_194 = _T_159 ? 5'h1c : _T_193; // @[Mux.scala 31:69:@153.4]
  assign _T_195 = _T_158 ? 5'h1b : _T_194; // @[Mux.scala 31:69:@154.4]
  assign _T_196 = _T_157 ? 5'h1a : _T_195; // @[Mux.scala 31:69:@155.4]
  assign _T_197 = _T_156 ? 5'h19 : _T_196; // @[Mux.scala 31:69:@156.4]
  assign _T_198 = _T_155 ? 5'h18 : _T_197; // @[Mux.scala 31:69:@157.4]
  assign _T_199 = _T_154 ? 5'h17 : _T_198; // @[Mux.scala 31:69:@158.4]
  assign _T_200 = _T_153 ? 5'h16 : _T_199; // @[Mux.scala 31:69:@159.4]
  assign _T_201 = _T_152 ? 5'h15 : _T_200; // @[Mux.scala 31:69:@160.4]
  assign _T_202 = _T_151 ? 5'h14 : _T_201; // @[Mux.scala 31:69:@161.4]
  assign _T_203 = _T_150 ? 5'h13 : _T_202; // @[Mux.scala 31:69:@162.4]
  assign _T_204 = _T_149 ? 5'h12 : _T_203; // @[Mux.scala 31:69:@163.4]
  assign _T_205 = _T_148 ? 5'h11 : _T_204; // @[Mux.scala 31:69:@164.4]
  assign _T_206 = _T_147 ? 5'h10 : _T_205; // @[Mux.scala 31:69:@165.4]
  assign _T_207 = _T_146 ? 5'hf : _T_206; // @[Mux.scala 31:69:@166.4]
  assign _T_208 = _T_145 ? 5'he : _T_207; // @[Mux.scala 31:69:@167.4]
  assign _T_209 = _T_144 ? 5'hd : _T_208; // @[Mux.scala 31:69:@168.4]
  assign _T_210 = _T_143 ? 5'hc : _T_209; // @[Mux.scala 31:69:@169.4]
  assign _T_211 = _T_142 ? 5'hb : _T_210; // @[Mux.scala 31:69:@170.4]
  assign _T_212 = _T_141 ? 5'ha : _T_211; // @[Mux.scala 31:69:@171.4]
  assign _T_213 = _T_140 ? 5'h9 : _T_212; // @[Mux.scala 31:69:@172.4]
  assign _T_214 = _T_139 ? 5'h8 : _T_213; // @[Mux.scala 31:69:@173.4]
  assign _T_215 = _T_138 ? 5'h7 : _T_214; // @[Mux.scala 31:69:@174.4]
  assign _T_216 = _T_137 ? 5'h6 : _T_215; // @[Mux.scala 31:69:@175.4]
  assign _T_217 = _T_136 ? 5'h5 : _T_216; // @[Mux.scala 31:69:@176.4]
  assign _T_218 = _T_135 ? 5'h4 : _T_217; // @[Mux.scala 31:69:@177.4]
  assign _T_219 = _T_134 ? 5'h3 : _T_218; // @[Mux.scala 31:69:@178.4]
  assign _T_220 = _T_133 ? 5'h2 : _T_219; // @[Mux.scala 31:69:@179.4]
  assign _T_221 = _T_132 ? 5'h1 : _T_220; // @[Mux.scala 31:69:@180.4]
  assign _T_222 = _T_131 ? 5'h0 : _T_221; // @[Mux.scala 31:69:@181.4]
  assign _T_223 = bits_to_decode[15:0]; // @[Bitwise.scala 109:18:@182.4]
  assign _T_228 = _T_223[15:8]; // @[Bitwise.scala 103:21:@185.4]
  assign _T_229 = {{8'd0}, _T_228}; // @[Bitwise.scala 103:31:@186.4]
  assign _T_230 = _T_223[7:0]; // @[Bitwise.scala 103:46:@187.4]
  assign _GEN_12 = {{8'd0}, _T_230}; // @[Bitwise.scala 103:65:@188.4]
  assign _T_231 = _GEN_12 << 8; // @[Bitwise.scala 103:65:@188.4]
  assign _T_233 = _T_231 & 16'hff00; // @[Bitwise.scala 103:75:@190.4]
  assign _T_234 = _T_229 | _T_233; // @[Bitwise.scala 103:39:@191.4]
  assign _T_238 = _T_234[15:4]; // @[Bitwise.scala 103:21:@195.4]
  assign _GEN_13 = {{4'd0}, _T_238}; // @[Bitwise.scala 103:31:@196.4]
  assign _T_239 = _GEN_13 & 16'hf0f; // @[Bitwise.scala 103:31:@196.4]
  assign _T_240 = _T_234[11:0]; // @[Bitwise.scala 103:46:@197.4]
  assign _GEN_14 = {{4'd0}, _T_240}; // @[Bitwise.scala 103:65:@198.4]
  assign _T_241 = _GEN_14 << 4; // @[Bitwise.scala 103:65:@198.4]
  assign _T_243 = _T_241 & 16'hf0f0; // @[Bitwise.scala 103:75:@200.4]
  assign _T_244 = _T_239 | _T_243; // @[Bitwise.scala 103:39:@201.4]
  assign _T_248 = _T_244[15:2]; // @[Bitwise.scala 103:21:@205.4]
  assign _GEN_15 = {{2'd0}, _T_248}; // @[Bitwise.scala 103:31:@206.4]
  assign _T_249 = _GEN_15 & 16'h3333; // @[Bitwise.scala 103:31:@206.4]
  assign _T_250 = _T_244[13:0]; // @[Bitwise.scala 103:46:@207.4]
  assign _GEN_16 = {{2'd0}, _T_250}; // @[Bitwise.scala 103:65:@208.4]
  assign _T_251 = _GEN_16 << 2; // @[Bitwise.scala 103:65:@208.4]
  assign _T_253 = _T_251 & 16'hcccc; // @[Bitwise.scala 103:75:@210.4]
  assign _T_254 = _T_249 | _T_253; // @[Bitwise.scala 103:39:@211.4]
  assign _T_258 = _T_254[15:1]; // @[Bitwise.scala 103:21:@215.4]
  assign _GEN_17 = {{1'd0}, _T_258}; // @[Bitwise.scala 103:31:@216.4]
  assign _T_259 = _GEN_17 & 16'h5555; // @[Bitwise.scala 103:31:@216.4]
  assign _T_260 = _T_254[14:0]; // @[Bitwise.scala 103:46:@217.4]
  assign _GEN_18 = {{1'd0}, _T_260}; // @[Bitwise.scala 103:65:@218.4]
  assign _T_261 = _GEN_18 << 1; // @[Bitwise.scala 103:65:@218.4]
  assign _T_263 = _T_261 & 16'haaaa; // @[Bitwise.scala 103:75:@220.4]
  assign _T_264 = _T_259 | _T_263; // @[Bitwise.scala 103:39:@221.4]
  assign _T_265 = bits_to_decode[30:16]; // @[Bitwise.scala 109:44:@222.4]
  assign _T_266 = _T_265[7:0]; // @[Bitwise.scala 109:18:@223.4]
  assign _T_271 = _T_266[7:4]; // @[Bitwise.scala 103:21:@226.4]
  assign _T_272 = {{4'd0}, _T_271}; // @[Bitwise.scala 103:31:@227.4]
  assign _T_273 = _T_266[3:0]; // @[Bitwise.scala 103:46:@228.4]
  assign _GEN_19 = {{4'd0}, _T_273}; // @[Bitwise.scala 103:65:@229.4]
  assign _T_274 = _GEN_19 << 4; // @[Bitwise.scala 103:65:@229.4]
  assign _T_276 = _T_274 & 8'hf0; // @[Bitwise.scala 103:75:@231.4]
  assign _T_277 = _T_272 | _T_276; // @[Bitwise.scala 103:39:@232.4]
  assign _T_281 = _T_277[7:2]; // @[Bitwise.scala 103:21:@236.4]
  assign _GEN_20 = {{2'd0}, _T_281}; // @[Bitwise.scala 103:31:@237.4]
  assign _T_282 = _GEN_20 & 8'h33; // @[Bitwise.scala 103:31:@237.4]
  assign _T_283 = _T_277[5:0]; // @[Bitwise.scala 103:46:@238.4]
  assign _GEN_21 = {{2'd0}, _T_283}; // @[Bitwise.scala 103:65:@239.4]
  assign _T_284 = _GEN_21 << 2; // @[Bitwise.scala 103:65:@239.4]
  assign _T_286 = _T_284 & 8'hcc; // @[Bitwise.scala 103:75:@241.4]
  assign _T_287 = _T_282 | _T_286; // @[Bitwise.scala 103:39:@242.4]
  assign _T_291 = _T_287[7:1]; // @[Bitwise.scala 103:21:@246.4]
  assign _GEN_22 = {{1'd0}, _T_291}; // @[Bitwise.scala 103:31:@247.4]
  assign _T_292 = _GEN_22 & 8'h55; // @[Bitwise.scala 103:31:@247.4]
  assign _T_293 = _T_287[6:0]; // @[Bitwise.scala 103:46:@248.4]
  assign _GEN_23 = {{1'd0}, _T_293}; // @[Bitwise.scala 103:65:@249.4]
  assign _T_294 = _GEN_23 << 1; // @[Bitwise.scala 103:65:@249.4]
  assign _T_296 = _T_294 & 8'haa; // @[Bitwise.scala 103:75:@251.4]
  assign _T_297 = _T_292 | _T_296; // @[Bitwise.scala 103:39:@252.4]
  assign _T_298 = _T_265[14:8]; // @[Bitwise.scala 109:44:@253.4]
  assign _T_299 = _T_298[3:0]; // @[Bitwise.scala 109:18:@254.4]
  assign _T_300 = _T_299[1:0]; // @[Bitwise.scala 109:18:@255.4]
  assign _T_301 = _T_300[0]; // @[Bitwise.scala 109:18:@256.4]
  assign _T_302 = _T_300[1]; // @[Bitwise.scala 109:44:@257.4]
  assign _T_304 = _T_299[3:2]; // @[Bitwise.scala 109:44:@259.4]
  assign _T_305 = _T_304[0]; // @[Bitwise.scala 109:18:@260.4]
  assign _T_306 = _T_304[1]; // @[Bitwise.scala 109:44:@261.4]
  assign _T_309 = _T_298[6:4]; // @[Bitwise.scala 109:44:@264.4]
  assign _T_310 = _T_309[1:0]; // @[Bitwise.scala 109:18:@265.4]
  assign _T_311 = _T_310[0]; // @[Bitwise.scala 109:18:@266.4]
  assign _T_312 = _T_310[1]; // @[Bitwise.scala 109:44:@267.4]
  assign _T_314 = _T_309[2]; // @[Bitwise.scala 109:44:@269.4]
  assign _T_318 = {_T_264,_T_297,_T_301,_T_302,_T_305,_T_306,_T_311,_T_312,_T_314}; // @[Cat.scala 30:58:@273.4]
  assign _T_319 = _T_318[0]; // @[OneHot.scala 39:40:@274.4]
  assign _T_320 = _T_318[1]; // @[OneHot.scala 39:40:@275.4]
  assign _T_321 = _T_318[2]; // @[OneHot.scala 39:40:@276.4]
  assign _T_322 = _T_318[3]; // @[OneHot.scala 39:40:@277.4]
  assign _T_323 = _T_318[4]; // @[OneHot.scala 39:40:@278.4]
  assign _T_324 = _T_318[5]; // @[OneHot.scala 39:40:@279.4]
  assign _T_325 = _T_318[6]; // @[OneHot.scala 39:40:@280.4]
  assign _T_326 = _T_318[7]; // @[OneHot.scala 39:40:@281.4]
  assign _T_327 = _T_318[8]; // @[OneHot.scala 39:40:@282.4]
  assign _T_328 = _T_318[9]; // @[OneHot.scala 39:40:@283.4]
  assign _T_329 = _T_318[10]; // @[OneHot.scala 39:40:@284.4]
  assign _T_330 = _T_318[11]; // @[OneHot.scala 39:40:@285.4]
  assign _T_331 = _T_318[12]; // @[OneHot.scala 39:40:@286.4]
  assign _T_332 = _T_318[13]; // @[OneHot.scala 39:40:@287.4]
  assign _T_333 = _T_318[14]; // @[OneHot.scala 39:40:@288.4]
  assign _T_334 = _T_318[15]; // @[OneHot.scala 39:40:@289.4]
  assign _T_335 = _T_318[16]; // @[OneHot.scala 39:40:@290.4]
  assign _T_336 = _T_318[17]; // @[OneHot.scala 39:40:@291.4]
  assign _T_337 = _T_318[18]; // @[OneHot.scala 39:40:@292.4]
  assign _T_338 = _T_318[19]; // @[OneHot.scala 39:40:@293.4]
  assign _T_339 = _T_318[20]; // @[OneHot.scala 39:40:@294.4]
  assign _T_340 = _T_318[21]; // @[OneHot.scala 39:40:@295.4]
  assign _T_341 = _T_318[22]; // @[OneHot.scala 39:40:@296.4]
  assign _T_342 = _T_318[23]; // @[OneHot.scala 39:40:@297.4]
  assign _T_343 = _T_318[24]; // @[OneHot.scala 39:40:@298.4]
  assign _T_344 = _T_318[25]; // @[OneHot.scala 39:40:@299.4]
  assign _T_345 = _T_318[26]; // @[OneHot.scala 39:40:@300.4]
  assign _T_346 = _T_318[27]; // @[OneHot.scala 39:40:@301.4]
  assign _T_347 = _T_318[28]; // @[OneHot.scala 39:40:@302.4]
  assign _T_348 = _T_318[29]; // @[OneHot.scala 39:40:@303.4]
  assign _T_381 = _T_348 ? 5'h1d : 5'h1e; // @[Mux.scala 31:69:@305.4]
  assign _T_382 = _T_347 ? 5'h1c : _T_381; // @[Mux.scala 31:69:@306.4]
  assign _T_383 = _T_346 ? 5'h1b : _T_382; // @[Mux.scala 31:69:@307.4]
  assign _T_384 = _T_345 ? 5'h1a : _T_383; // @[Mux.scala 31:69:@308.4]
  assign _T_385 = _T_344 ? 5'h19 : _T_384; // @[Mux.scala 31:69:@309.4]
  assign _T_386 = _T_343 ? 5'h18 : _T_385; // @[Mux.scala 31:69:@310.4]
  assign _T_387 = _T_342 ? 5'h17 : _T_386; // @[Mux.scala 31:69:@311.4]
  assign _T_388 = _T_341 ? 5'h16 : _T_387; // @[Mux.scala 31:69:@312.4]
  assign _T_389 = _T_340 ? 5'h15 : _T_388; // @[Mux.scala 31:69:@313.4]
  assign _T_390 = _T_339 ? 5'h14 : _T_389; // @[Mux.scala 31:69:@314.4]
  assign _T_391 = _T_338 ? 5'h13 : _T_390; // @[Mux.scala 31:69:@315.4]
  assign _T_392 = _T_337 ? 5'h12 : _T_391; // @[Mux.scala 31:69:@316.4]
  assign _T_393 = _T_336 ? 5'h11 : _T_392; // @[Mux.scala 31:69:@317.4]
  assign _T_394 = _T_335 ? 5'h10 : _T_393; // @[Mux.scala 31:69:@318.4]
  assign _T_395 = _T_334 ? 5'hf : _T_394; // @[Mux.scala 31:69:@319.4]
  assign _T_396 = _T_333 ? 5'he : _T_395; // @[Mux.scala 31:69:@320.4]
  assign _T_397 = _T_332 ? 5'hd : _T_396; // @[Mux.scala 31:69:@321.4]
  assign _T_398 = _T_331 ? 5'hc : _T_397; // @[Mux.scala 31:69:@322.4]
  assign _T_399 = _T_330 ? 5'hb : _T_398; // @[Mux.scala 31:69:@323.4]
  assign _T_400 = _T_329 ? 5'ha : _T_399; // @[Mux.scala 31:69:@324.4]
  assign _T_401 = _T_328 ? 5'h9 : _T_400; // @[Mux.scala 31:69:@325.4]
  assign _T_402 = _T_327 ? 5'h8 : _T_401; // @[Mux.scala 31:69:@326.4]
  assign _T_403 = _T_326 ? 5'h7 : _T_402; // @[Mux.scala 31:69:@327.4]
  assign _T_404 = _T_325 ? 5'h6 : _T_403; // @[Mux.scala 31:69:@328.4]
  assign _T_405 = _T_324 ? 5'h5 : _T_404; // @[Mux.scala 31:69:@329.4]
  assign _T_406 = _T_323 ? 5'h4 : _T_405; // @[Mux.scala 31:69:@330.4]
  assign _T_407 = _T_322 ? 5'h3 : _T_406; // @[Mux.scala 31:69:@331.4]
  assign _T_408 = _T_321 ? 5'h2 : _T_407; // @[Mux.scala 31:69:@332.4]
  assign _T_409 = _T_320 ? 5'h1 : _T_408; // @[Mux.scala 31:69:@333.4]
  assign _T_410 = _T_319 ? 5'h0 : _T_409; // @[Mux.scala 31:69:@334.4]
  assign number_of_same_bit_value = _T_33 ? _T_222 : _T_410; // @[POSIT.scala 80:36:@335.4]
  assign _T_413 = bits_to_decode[0]; // @[POSIT.scala 98:47:@338.4]
  assign _T_417 = number_of_same_bit_value == 5'h1e; // @[POSIT.scala 98:84:@340.4]
  assign _T_418 = _T_413 & _T_417; // @[POSIT.scala 98:57:@341.4]
  assign _T_419 = {1'b0,$signed(number_of_same_bit_value)}; // @[POSIT.scala 99:58:@342.4]
  assign _T_422 = $signed(_T_419) - $signed(6'sh1); // @[POSIT.scala 100:63:@344.4]
  assign _T_423 = $signed(_T_419) - $signed(6'sh1); // @[POSIT.scala 100:63:@345.4]
  assign _T_424 = $signed(_T_423); // @[POSIT.scala 100:63:@346.4]
  assign _T_425 = _T_418 ? $signed(_T_419) : $signed(_T_424); // @[POSIT.scala 98:32:@347.4]
  assign _T_428 = _T_413 == 1'h0; // @[POSIT.scala 101:51:@349.4]
  assign _T_431 = _T_428 & _T_417; // @[POSIT.scala 101:58:@351.4]
  assign _T_434 = $signed(6'sh0) - $signed(_T_419); // @[POSIT.scala 102:30:@353.4]
  assign _T_435 = $signed(6'sh0) - $signed(_T_419); // @[POSIT.scala 102:30:@354.4]
  assign _T_436 = $signed(_T_435); // @[POSIT.scala 102:30:@355.4]
  assign _T_438 = $signed(_T_436) - $signed(6'sh1); // @[POSIT.scala 102:61:@356.4]
  assign _T_439 = $signed(_T_436) - $signed(6'sh1); // @[POSIT.scala 102:61:@357.4]
  assign _T_440 = $signed(_T_439); // @[POSIT.scala 102:61:@358.4]
  assign _T_446 = _T_431 ? $signed(_T_440) : $signed(_T_436); // @[POSIT.scala 101:33:@363.4]
  assign _T_447 = _T_33 ? $signed(_T_425) : $signed(_T_446); // @[POSIT.scala 97:29:@364.4]
  assign _T_449 = number_of_same_bit_value + 5'h1; // @[POSIT.scala 108:56:@366.4]
  assign _T_454 = $signed(7'sh20) - $signed(7'sh1); // @[POSIT.scala 116:37:@370.4]
  assign _T_455 = $signed(7'sh20) - $signed(7'sh1); // @[POSIT.scala 116:37:@371.4]
  assign _T_456 = $signed(_T_455); // @[POSIT.scala 116:37:@372.4]
  assign _T_457 = {1'b0,$signed(io_o_posit_regime_size)}; // @[POSIT.scala 116:68:@373.4]
  assign _GEN_24 = {{1{_T_457[5]}},_T_457}; // @[POSIT.scala 116:43:@374.4]
  assign _T_458 = $signed(_T_456) - $signed(_GEN_24); // @[POSIT.scala 116:43:@374.4]
  assign _T_459 = $signed(_T_456) - $signed(_GEN_24); // @[POSIT.scala 116:43:@375.4]
  assign _T_460 = $signed(_T_459); // @[POSIT.scala 116:43:@376.4]
  assign _T_461 = {1'b0,$signed(io_o_posit_max_exponent_size)}; // @[POSIT.scala 116:104:@377.4]
  assign _GEN_25 = {{1{_T_461[5]}},_T_461}; // @[POSIT.scala 116:73:@378.4]
  assign _T_462 = $signed(_T_460) - $signed(_GEN_25); // @[POSIT.scala 116:73:@378.4]
  assign _T_463 = $signed(_T_460) - $signed(_GEN_25); // @[POSIT.scala 116:73:@379.4]
  assign _T_464 = $signed(_T_463); // @[POSIT.scala 116:73:@380.4]
  assign _GEN_26 = _T_464[5:0]; // @[POSIT.scala 115:37:@369.4 POSIT.scala 116:27:@381.4]
  assign posible_fraction_size = $signed(_GEN_26); // @[POSIT.scala 115:37:@369.4 POSIT.scala 116:27:@381.4]
  assign _T_466 = $signed(posible_fraction_size) <= $signed(6'sh0); // @[POSIT.scala 117:59:@382.4]
  assign _T_470 = 6'h20 - 6'h1; // @[POSIT.scala 119:44:@383.4]
  assign _T_471 = $unsigned(_T_470); // @[POSIT.scala 119:44:@384.4]
  assign _T_472 = _T_471[5:0]; // @[POSIT.scala 119:44:@385.4]
  assign _GEN_27 = {{1'd0}, io_o_posit_regime_size}; // @[POSIT.scala 119:50:@386.4]
  assign _T_473 = _T_472 - _GEN_27; // @[POSIT.scala 119:50:@386.4]
  assign _T_474 = $unsigned(_T_473); // @[POSIT.scala 119:50:@387.4]
  assign _T_475 = _T_474[5:0]; // @[POSIT.scala 119:50:@388.4]
  assign _GEN_28 = {{1'd0}, io_o_posit_max_exponent_size}; // @[POSIT.scala 119:75:@389.4]
  assign _T_476 = _T_475 - _GEN_28; // @[POSIT.scala 119:75:@389.4]
  assign _T_477 = $unsigned(_T_476); // @[POSIT.scala 119:75:@390.4]
  assign _T_478 = _T_477[5:0]; // @[POSIT.scala 119:75:@391.4]
  assign _T_479 = _T_466 ? 6'h0 : _T_478; // @[POSIT.scala 117:36:@392.4]
  assign _T_481 = io_o_posit_fraction_size == 5'h0; // @[POSIT.scala 124:57:@394.4]
  assign _GEN_29 = {{1'd0}, io_o_posit_fraction_size}; // @[POSIT.scala 126:65:@396.4]
  assign _T_489 = 6'h20 - _GEN_29; // @[POSIT.scala 126:65:@396.4]
  assign _T_490 = $unsigned(_T_489); // @[POSIT.scala 126:65:@397.4]
  assign _T_491 = _T_490[5:0]; // @[POSIT.scala 126:65:@398.4]
  assign _T_492 = 32'hffffffff >> _T_491; // @[POSIT.scala 126:55:@399.4]
  assign _GEN_30 = {{1'd0}, bits_to_decode}; // @[POSIT.scala 126:92:@400.4]
  assign _T_493 = _T_492 & _GEN_30; // @[POSIT.scala 126:92:@400.4]
  assign _GEN_32 = _T_460[5:0]; // @[POSIT.scala 131:39:@403.4 POSIT.scala 132:29:@411.4]
  assign posible_exponent_size_1 = $signed(_GEN_32); // @[POSIT.scala 131:39:@403.4 POSIT.scala 132:29:@411.4]
  assign _T_507 = $signed(posible_exponent_size_1) < $signed(_T_461); // @[POSIT.scala 134:60:@414.4]
  assign posible_exponent_size_2 = _T_507 ? $signed(posible_exponent_size_1) : $signed(_T_461); // @[POSIT.scala 134:35:@416.4]
  assign _T_511 = $signed(posible_exponent_size_2) <= $signed(6'sh0); // @[POSIT.scala 137:61:@418.4]
  assign _T_513 = $unsigned(posible_exponent_size_2); // @[POSIT.scala 139:61:@419.4]
  assign _T_514 = _T_511 ? 6'h0 : _T_513; // @[POSIT.scala 137:36:@420.4]
  assign _T_516 = io_o_posit_exponent_size == 5'h0; // @[POSIT.scala 146:57:@422.4]
  assign _T_518 = bits_to_decode >> io_o_posit_fraction_size; // @[POSIT.scala 148:48:@423.4]
  assign _GEN_33 = {{1'd0}, io_o_posit_exponent_size}; // @[POSIT.scala 149:64:@425.4]
  assign _T_525 = 6'h20 - _GEN_33; // @[POSIT.scala 149:64:@425.4]
  assign _T_526 = $unsigned(_T_525); // @[POSIT.scala 149:64:@426.4]
  assign _T_527 = _T_526[5:0]; // @[POSIT.scala 149:64:@427.4]
  assign _T_528 = 32'hffffffff >> _T_527; // @[POSIT.scala 149:53:@428.4]
  assign _GEN_34 = {{1'd0}, _T_518}; // @[POSIT.scala 148:79:@429.4]
  assign _T_529 = _GEN_34 & _T_528; // @[POSIT.scala 148:79:@429.4]
  assign io_o_posit_sign = io_i_bits[31]; // @[POSIT.scala 54:21:@16.4]
  assign io_o_posit_special_number = _T_14 | _T_17; // @[POSIT.scala 47:31:@14.4]
  assign io_o_posit_regime = {{26{_T_447[5]}},_T_447}; // @[POSIT.scala 97:23:@365.4]
  assign io_o_posit_exponent = _T_516 ? 32'h0 : _T_529; // @[POSIT.scala 146:25:@431.4]
  assign io_o_posit_fraction = _T_481 ? 32'h0 : _T_493; // @[POSIT.scala 124:25:@402.4]
  assign io_o_posit_regime_size = number_of_same_bit_value + 5'h1; // @[POSIT.scala 108:28:@368.4]
  assign io_o_posit_exponent_size = _T_514[4:0]; // @[POSIT.scala 137:30:@421.4]
  assign io_o_posit_fraction_size = _T_479[4:0]; // @[POSIT.scala 117:30:@393.4]
  assign io_o_posit_max_exponent_size = 5'h3; // @[POSIT.scala 63:34:@18.4]
endmodule
